 
module transform ();

endmodule