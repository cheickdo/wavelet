module mult(
    input [size-1:0] in0,
    input [size-1:0] in1,
    output [size-1:0] product
);
    

endmodule