
//cumulative pipelined adder
module cummadd();

endmodule