
//Divider module
module div(
    input [size-1::0] in,
    output reg [size-1::0] out
);

    parameter size = 32;
    
    //

endmodule